module Instr_mem(input logic [31:0] a,
					output logic [31:0] rd);

reg [31:0] RAM [23:0];
logic [31:0] data;

assign rd = data;

initial
	$readmemh("memfile.dat",RAM);

always_ff @(a)
begin : MEM_READ
	data <= RAM[a[31:2]];
end

endmodule 